library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC.STD.ALL;

entity RAM is
  port(
    Clk   :in STD_LOGIC;
    Rst   :in STD_LOGIC;
    EN    :in STD_LOGIC;
    x     :in STD_LOGIC_VECTOR(15 downto 0);
    y     :out STD_LOGIC_VECTOR(15 downto 0)
  );
 end entity;
    
 architecture behavioral of RAM is
 end behavioral;
