library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC.STD.ALL;

entity RAM is
  port(
    );
 end entity;
    
 architecture behavioral of RAM is
 end behavioral;
